module color_map (
    input [7:0] color,
    output [23:0] rgb
);
    
endmodule